module mux (sel, res);
	input  [2:0] sel;
	output [7:0] res;
	reg    [7:0] res;
	always @(sel or res) begin
	   case (sel)
	      3’b000  : res = 8’b00000001;
	      3’b001  : res = 8’b00000010;
	      3’b010  : res = 8’b00000100;
	      3’b011  : res = 8’b00001000;
	      3’b100  : res = 8’b00010000;
	      3’b101  : res = 8’b00100000;
	      // 110 and 111 selector values are unused
	      default : res = 8’bxxxxxxxx;
	   endcase
	end
        endmodule
